module and_R (
				input logic A,B,
				output logic y
				);
				
assign y = A & B;
endmodule
				